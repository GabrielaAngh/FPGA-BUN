library verilog;
use verilog.vl_types.all;
entity test_sync is
end test_sync;
